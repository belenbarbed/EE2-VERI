module fsm (
		clk,
		tick,
		trigger,
		time_out,
		en_lfsr,
		start_delay,
		ledr
);

	input clk;
	input tick;
	input trigger;
	input time_out;
	
	output en_lfsr;
	output start_delay;
	output [9:0] ledr;
	
	




endmodule 