module delay (
		N,
		clk,
		trigger,
		time_out
);

	input [6:0] N;
	input clk;
	input trigger;
	
	output time_out;



endmodule 